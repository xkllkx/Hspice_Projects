**Trans_OR**
.subckt  T_OR  input1  input2  output  wmin

MP1  node1   input1  vdd     vdd   pmos  l=90n    w=3*wmin
MN1  node1   input1  gnd     gnd   nmos  l=90n    w=wmin

MP2  output  input1  input2  vdd   pmos  l=90n    w=3*wmin
MN2  input2  node1   output  gnd   nmos  l=90n    w=wmin

MP3  output  node1   input1  vdd   pmos  l=90n    w=3*wmin

.ends
